netcdf MTP {
dimensions:
	MTPTime = UNLIMITED ; 
	Time = UNLIMITED ; 
	MTPTpl = 30 ;		/// the number of templates created for the MTP
	ALT_MTP = 33 ;		/// the Altitude coordinate variable for profiles
	TPLALT_MTP = 33;	/// the flight level Altitudes for templates
	TPLIDX_MTP = 43;	/// index into templates
	MTPChan = 3 ;		/// the number of frequency channels for the MTP
	BTSCANANGLE_MTP = 10 ;	/// for Brightness Temperatures
	CNTSCANANGLE_MTP = 12 ;	/// for Raw Scans including 2 target counts
variables:
	int MTPTime(MTPTime) ;
		MTPTime:long_name = "time of MTP measurement" ;
		MTPTime:standard_name = "time" ;
		MTPTime:units = "seconds since 2014-07-20 00:00:00 +0000" ;
		MTPTime:strptime_format = "seconds since %F %T %z" ;
	int Time(Time) ;
		Time:long_name = "time of measurement" ;
		Time:standard_name = "time" ;
		Time:units = "seconds since 2014-07-20 00:00:00 +0000" ;
		Time:strptime_format = "seconds since %F %T %z" ;
	float CNTSCANANGLE_MTP(CNTSCANANGLE_MTP) ;
		CNTSCANANGLE_MTP:long_name = "MTP Pointing Angle (incl Target)" ;
		CNTSCANANGLE_MTP:units = "degree" ;
		CNTSCANANGLE_MTP:valid_range = -180.f, 90.f ;
	float CNT_MTP(MTPTime, MTPChan, CNTSCANANGLE_MTP) ;
		CNT_MTP:_FillValue = -32767.f ;
		CNT_MTP:units = "count" ;
		CNT_MTP:long_name = "MTP Channel Scan Counts (incl Target)" ;
		CNT_MTP:Category = "MTP" ;
	float BTSCANANGLE_MTP(BTSCANANGLE_MTP) ; 
		BTSCANANGLE_MTP:long_name = "MTP Pointing Angle" ;
		BTSCANANGLE_MTP:units = "degree" ;
		BTSCANANGLE_MTP:valid_range = -90.f, 90.f ;
	float BT_MTP(MTPTime, MTPChan, BTSCANANGLE_MTP) ;
		BT_MTP:_FillValue = -32767.f ;
		BT_MTP:units = "deg_K" ;
		BT_MTP:long_name = "MTP Brightness Temperatures" ;
		BT_MTP:Category = "MTP" ;
	int TPLIDX_MTP(MTPTime) ;    // Primary template index used to generate this profile
	int TPLIDX2_MTP(MTPTime) ;   // 2ndary template index (if used) to generate this profile
		TPLIDX2_MTP:_FillValue = -32767 ; // Indicates not used
	float TPLALT_MTP(MTPTime, TPLALT_MTP) ;   // Template Altitude used
		TPLALT_MTP:long_name = "MTP Template Altitude" ;
		TPLALT_MTP:units = "km" ;
	float TPLBT_MTP(TPLIDX_MTP, TPLALT_MTP, MTPChan, BTSCANANGLE_MTP) ;
		TPLBT_MTP:_FillValue = -32767.f ;
		TPLBT_MTP:units = "deg_K" ;
		TPLBT_MTP:long_name = "MTP Template Brightness Temperature" ;
		TPLBT_MTP:Category = "MTP" ;
        string TPLID_MTP(TPLIDX_MTP) ;  // Template identifier
	string TPLOBSTIME_MTP(MTPTpl) ;
		TPLOBSTIME_MTP:units = "ISO 8601 UTC string" ;
	float TPLLAT_MTP(MTPTpl) ;
		TPLLAT_MTP:_FillValue = -32767.f ;
		TPLLAT_MTP:units = "degree_N" ;
		TPLLAT_MTP:long_name = "Latitude of Rawindsonde used for template" ;
	float TPLLON_MTP(MTPTpl) ;
		TPLLON_MTP:_FillValue = -32767.f ;
		TPLLON_MTP:units = "degree_E" ;
		TPLLON_MTP:long_name = "Longitude of Rawindsonde used for template" ;
	float ALT_MTP(MTPTime, ALT_MTP) ;
		ALT_MTP:_FillValue = -32767.f ;
		ALT_MTP:units = "km" ;
		ALT_MTP:long_name = "MTP ATP Altitude" ;
		ALT_MTP:standard_name = "altitude" ;
		ALT_MTP:Category = "MTP" ;
	float TEMP_MTP(MTPTime, ALT_MTP) ;
		TEMP_MTP:_FillValue = -32767.f ;
		TEMP_MTP:units = "deg_K" ;
		TEMP_MTP:long_name = "MTP ATP Temperature" ;
		TEMP_MTP:Category = "MTP" ;
	float MRI_MTP(MTPTime) ;
		MRI_MTP:_FillValue = -32767.f ;
		MRI_MTP:units = "count" ;
		MRI_MTP:long_name = "MTP Quality Indicator" ;
		MRI_MTP:actual_range = 0.f, 2.f ;
		MRI_MTP:Category = "MTP" ;
	float MTPFREQ(MTPChan) ;
		MTPFREQ:units = "GHz";
	float ACCPCNTE_MTP(MTPTime) ;
		ACCPCNTE_MTP:_FillValue = -32767.f ;
		ACCPCNTE_MTP:units = "count" ;
		ACCPCNTE_MTP:long_name = "MTP Engineering Multiplxr Acceler Counts" ;
		ACCPCNTE_MTP:actual_range = 1548.f, 2238.f ;
		ACCPCNTE_MTP:Category = "MTP" ;
	float SMCMD_MTP(MTPTime) ;
		SMCMD_MTP:_FillValue = -32767.f ;
		SMCMD_MTP:units = "count" ;
		SMCMD_MTP:long_name = "MTP Scan Motor Commanded Position" ;
		SMCMD_MTP:actual_range = 72196.f, 79364.f ;
		SMCMD_MTP:Category = "MTP" ;
	float SMENC_MTP(MTPTime) ;
		SMENC_MTP:_FillValue = -32767.f ;
		SMENC_MTP:units = "count" ;
		SMENC_MTP:long_name = "MTP Scan Motor Encoded Position" ;
		SMENC_MTP:actual_range = 71232.f, 78864.f ;
		SMENC_MTP:Category = "MTP" ;
	float TAIRCNTE_MTP(MTPTime) ;
		TAIRCNTE_MTP:_FillValue = -32767.f ;
		TAIRCNTE_MTP:units = "count" ;
		TAIRCNTE_MTP:long_name = "MTP Engineering Multiplxr T Pod Air Counts" ;
		TAIRCNTE_MTP:actual_range = 2461.f, 3077.f ;
		TAIRCNTE_MTP:Category = "MTP" ;
	float TAMPCNTP_MTP(MTPTime) ;
		TAMPCNTP_MTP:_FillValue = -32767.f ;
		TAMPCNTP_MTP:units = "count" ;
		TAMPCNTP_MTP:long_name = "MTP Platinum Multiplxr Amplifier Temp Counts" ;
		TAMPCNTP_MTP:actual_range = 13292.f, 13488.f ;
		TAMPCNTP_MTP:Category = "MTP" ;
	float TDATCNTE_MTP(MTPTime) ;
		TDATCNTE_MTP:_FillValue = -32767.f ;
		TDATCNTE_MTP:units = "count" ;
		TDATCNTE_MTP:long_name = "MTP Engineering Multiplxr T Data Counts" ;
		TDATCNTE_MTP:actual_range = 1282.f, 1424.f ;
		TDATCNTE_MTP:Category = "MTP" ;
	float TMIXCNTP_MTP(MTPTime) ;
		TMIXCNTP_MTP:_FillValue = -32767.f ;
		TMIXCNTP_MTP:units = "count" ;
		TMIXCNTP_MTP:long_name = "MTP Platinum Multiplxr Mixer Temperature Counts" ;
		TMIXCNTP_MTP:actual_range = 13312.f, 13497.f ;
		TMIXCNTP_MTP:Category = "MTP" ;
	float TMTRCNTE_MTP(MTPTime) ;
		TMTRCNTE_MTP:_FillValue = -32767.f ;
		TMTRCNTE_MTP:units = "count" ;
		TMTRCNTE_MTP:long_name = "MTP Engineering Multiplxr T Motor Counts" ;
		TMTRCNTE_MTP:actual_range = 2312.f, 2809.f ;
		TMTRCNTE_MTP:Category = "MTP" ;
	float TNCCNTE_MTP(MTPTime) ;
		TNCCNTE_MTP:_FillValue = -32767.f ;
		TNCCNTE_MTP:units = "count" ;
		TNCCNTE_MTP:long_name = "MTP Engineering Multiplxr T N/C Counts" ;
		TNCCNTE_MTP:actual_range = 4095.f, 4095.f ;
		TNCCNTE_MTP:Category = "MTP" ;
	float TNDCNTP_MTP(MTPTime) ;
		TNDCNTP_MTP:_FillValue = -32767.f ;
		TNDCNTP_MTP:units = "count" ;
		TNDCNTP_MTP:long_name = "MTP Platinum Multiplxr Noise Diode Temp Counts" ;
		TNDCNTP_MTP:actual_range = 13095.f, 13308.f ;
		TNDCNTP_MTP:Category = "MTP" ;
	float TPSPCNTE_MTP(MTPTime) ;
		TPSPCNTE_MTP:_FillValue = -32767.f ;
		TPSPCNTE_MTP:units = "count" ;
		TPSPCNTE_MTP:long_name = "MTP Engineering Multiplxr T Power Supply Counts" ;
		TPSPCNTE_MTP:actual_range = 1541.f, 1677.f ;
		TPSPCNTE_MTP:Category = "MTP" ;
	float TR350CNTP_MTP(MTPTime) ;
		TR350CNTP_MTP:_FillValue = -32767.f ;
		TR350CNTP_MTP:units = "count" ;
		TR350CNTP_MTP:long_name = "MTP Platinum Multiplxr R350 Counts" ;
		TR350CNTP_MTP:actual_range = 2165.f, 2176.f ;
		TR350CNTP_MTP:Category = "MTP" ;
	float TR600CNTP_MTP(MTPTime) ;
		TR600CNTP_MTP:_FillValue = -32767.f ;
		TR600CNTP_MTP:units = "count" ;
		TR600CNTP_MTP:long_name = "MTP Platinum Multiplxr R600 Counts" ;
		TR600CNTP_MTP:actual_range = 14442.f, 14463.f ;
		TR600CNTP_MTP:Category = "MTP" ;
	float TSMPCNTE_MTP(MTPTime) ;
		TSMPCNTE_MTP:_FillValue = -32767.f ;
		TSMPCNTE_MTP:units = "count" ;
		TSMPCNTE_MTP:long_name = "MTP Engineering Multiplxr T Scan Counts" ;
		TSMPCNTE_MTP:actual_range = 2469.f, 3145.f ;
		TSMPCNTE_MTP:Category = "MTP" ;
	float TSYNCNTE_MTP(MTPTime) ;
		TSYNCNTE_MTP:_FillValue = -32767.f ;
		TSYNCNTE_MTP:units = "count" ;
		TSYNCNTE_MTP:long_name = "MTP Engineering Multiplxr T Synth Counts" ;
		TSYNCNTE_MTP:actual_range = 1511.f, 1621.f ;
		TSYNCNTE_MTP:Category = "MTP" ;
	float TTCNTRCNTP_MTP(MTPTime) ;
		TTCNTRCNTP_MTP:_FillValue = -32767.f ;
		TTCNTRCNTP_MTP:units = "count" ;
		TTCNTRCNTP_MTP:long_name = "MTP Platinum Multiplxr Target Center Temp Counts" ;
		TTCNTRCNTP_MTP:actual_range = 13793.f, 13823.f ;
		TTCNTRCNTP_MTP:Category = "MTP" ;
	float TTEDGCNTP_MTP(MTPTime) ;
		TTEDGCNTP_MTP:_FillValue = -32767.f ;
		TTEDGCNTP_MTP:units = "count" ;
		TTEDGCNTP_MTP:long_name = "MTP Platinum Multiplxr Target Edge Temp Counts" ;
		TTEDGCNTP_MTP:actual_range = 13784.f, 13817.f ;
		TTEDGCNTP_MTP:Category = "MTP" ;
	float TWINCNTP_MTP(MTPTime) ;
		TWINCNTP_MTP:_FillValue = -32767.f ;
		TWINCNTP_MTP:units = "count" ;
		TWINCNTP_MTP:long_name = "MTP Platinum Multiplxr Polyethelene Window Temp Counts" ;
		TWINCNTP_MTP:actual_range = 6788.f, 10190.f ;
		TWINCNTP_MTP:Category = "MTP" ;
	float VM08CNTE_MTP(MTPTime) ;
		VM08CNTE_MTP:_FillValue = -32767.f ;
		VM08CNTE_MTP:units = "count" ;
		VM08CNTE_MTP:long_name = "MTP Engineering Multiplxr Vm08 Counts" ;
		VM08CNTE_MTP:actual_range = 2927.f, 2928.f ;
		VM08CNTE_MTP:Category = "MTP" ;
	float VM15CNTE_MTP(MTPTime) ;
		VM15CNTE_MTP:_FillValue = -32767.f ;
		VM15CNTE_MTP:units = "count" ;
		VM15CNTE_MTP:long_name = "MTP Engineering Multiplxr VM15 Counts" ;
		VM15CNTE_MTP:actual_range = 2941.f, 2945.f ;
		VM15CNTE_MTP:Category = "MTP" ;
	float VMTRCNTE_MTP(MTPTime) ;
		VMTRCNTE_MTP:_FillValue = -32767.f ;
		VMTRCNTE_MTP:units = "count" ;
		VMTRCNTE_MTP:long_name = "MTP Engineering Multiplxr Vmtr Counts" ;
		VMTRCNTE_MTP:actual_range = 3075.f, 3091.f ;
		VMTRCNTE_MTP:Category = "MTP" ;
	float VP05CNTE_MTP(MTPTime) ;
		VP05CNTE_MTP:_FillValue = -32767.f ;
		VP05CNTE_MTP:units = "count" ;
		VP05CNTE_MTP:long_name = "MTP Engineering Multiplxr Vp05 Counts" ;
		VP05CNTE_MTP:actual_range = 2428.f, 2433.f ;
		VP05CNTE_MTP:Category = "MTP" ;
	float VP08CNTE_MTP(MTPTime) ;
		VP08CNTE_MTP:_FillValue = -32767.f ;
		VP08CNTE_MTP:units = "count" ;
		VP08CNTE_MTP:long_name = "MTP Engineering Multiplxr Vp08 Counts" ;
		VP08CNTE_MTP:actual_range = 2898.f, 2899.f ;
		VP08CNTE_MTP:Category = "MTP" ;
	float VP15CNTE_MTP(MTPTime) ;
		VP15CNTE_MTP:_FillValue = -32767.f ;
		VP15CNTE_MTP:units = "count" ;
		VP15CNTE_MTP:long_name = "MTP Engineering Multiplxr Vp15 Counts" ;
		VP15CNTE_MTP:actual_range = 2908.f, 2928.f ;
		VP15CNTE_MTP:Category = "MTP" ;
	float VSYNCNTE_MTP(MTPTime) ;
		VSYNCNTE_MTP:_FillValue = -32767.f ;
		VSYNCNTE_MTP:units = "count" ;
		VSYNCNTE_MTP:long_name = "MTP Engineering Multiplxr Vsyn Counts" ;
		VSYNCNTE_MTP:actual_range = 1920.f, 1932.f ;
		VSYNCNTE_MTP:Category = "MTP" ;
	float VVIDCNTE_MTP(MTPTime) ;
		VVIDCNTE_MTP:_FillValue = -32767.f ;
		VVIDCNTE_MTP:units = "count" ;
		VVIDCNTE_MTP:long_name = "MTP Engineering Multiplxr Vvid Counts" ;
		VVIDCNTE_MTP:actual_range = 2084.f, 2352.f ;
		VVIDCNTE_MTP:Category = "MTP" ;
///  The following are probably unnecessary.  They are currently coming from the Visual Basic
///  UDP feed.  They could be nice to have for comparison w/VB MTP
	float PDAY_MTP(MTPTime) ;
		PDAY_MTP:_FillValue = -32767.f ;
		PDAY_MTP:units = "count" ;
		PDAY_MTP:long_name = "MTP ATP Day" ;
		PDAY_MTP:actual_range = 20.f, 20.f ;
		PDAY_MTP:Category = "MTP" ;
	float PHOUR_MTP(MTPTime) ;
		PHOUR_MTP:_FillValue = -32767.f ;
		PHOUR_MTP:units = "count" ;
		PHOUR_MTP:long_name = "MTP ATP Hour" ;
		PHOUR_MTP:actual_range = 8.f, 14.f ;
		PHOUR_MTP:Category = "MTP" ;
	float PMIN_MTP(MTPTime) ;
		PMIN_MTP:_FillValue = -32767.f ;
		PMIN_MTP:units = "count" ;
		PMIN_MTP:long_name = "MTP ATP Minute" ;
		PMIN_MTP:actual_range = 0.f, 59.f ;
		PMIN_MTP:Category = "MTP" ;
	float PMONTH_MTP(MTPTime) ;
		PMONTH_MTP:_FillValue = -32767.f ;
		PMONTH_MTP:units = "count" ;
		PMONTH_MTP:long_name = "MTP ATP Month" ;
		PMONTH_MTP:actual_range = 7.f, 7.f ;
		PMONTH_MTP:Category = "MTP" ;
	float PSEC_MTP(MTPTime) ;
		PSEC_MTP:_FillValue = -32767.f ;
		PSEC_MTP:units = "count" ;
		PSEC_MTP:long_name = "MTP ATP Second" ;
		PSEC_MTP:actual_range = 0.f, 59.f ;
		PSEC_MTP:Category = "MTP" ;
	float PYEAR_MTP(MTPTime) ;
		PYEAR_MTP:_FillValue = -32767.f ;
		PYEAR_MTP:units = "count" ;
		PYEAR_MTP:long_name = "MTP ATP Year" ;
		PYEAR_MTP:actual_range = 2014.f, 2014.f ;
		PYEAR_MTP:Category = "MTP" ;
	float SAAT_MTP(MTPTime) ;
		SAAT_MTP:_FillValue = -32767.f ;
		SAAT_MTP:units = "deg_K" ;
		SAAT_MTP:long_name = "MTP Scan Avg Ambient Air Temp" ;
		SAAT_MTP:actual_range = 218.08f, 278.5f ;
		SAAT_MTP:Category = "MTP" ;
	float SALAT_MTP(MTPTime) ;
		SALAT_MTP:_FillValue = -32767.f ;
		SALAT_MTP:units = "degree_N" ;
		SALAT_MTP:long_name = "MTP Scan Avg Latitude" ;
		SALAT_MTP:actual_range = -46.32f, -41.86f ;
		SALAT_MTP:Category = "MTP" ;
	float SALON_MTP(MTPTime) ;
		SALON_MTP:_FillValue = -32767.f ;
		SALON_MTP:units = "degree_E" ;
		SALON_MTP:long_name = "MTP Scan Avg Longitude" ;
		SALON_MTP:actual_range = 165.219f, 173.261f ;
		SALON_MTP:Category = "MTP" ;
	float SAPALT_MTP(MTPTime) ;
		SAPALT_MTP:_FillValue = -32767.f ;
		SAPALT_MTP:units = "km" ;
		SAPALT_MTP:long_name = "MTP Scan Avg Pressure Altitude" ;
		SAPALT_MTP:actual_range = 0.09f, 12.19f ;
		SAPALT_MTP:Category = "MTP" ;
	float SAPITCH_MTP(MTPTime) ;
		SAPITCH_MTP:_FillValue = -32767.f ;
		SAPITCH_MTP:units = "degree" ;
		SAPITCH_MTP:long_name = "MTP Scan Avg Pitch" ;
		SAPITCH_MTP:actual_range = -2.33f, 14.52f ;
		SAPITCH_MTP:Category = "MTP" ;
	float SAROLL_MTP(MTPTime) ;
		SAROLL_MTP:_FillValue = -32767.f ;
		SAROLL_MTP:units = "degree" ;
		SAROLL_MTP:long_name = "MTP Scan Avg Roll" ;
		SAROLL_MTP:actual_range = -22.99f, 25.28f ;
		SAROLL_MTP:Category = "MTP" ;
	float SDAY_MTP(MTPTime) ;
		SDAY_MTP:_FillValue = -32767.f ;
		SDAY_MTP:units = "count" ;
		SDAY_MTP:long_name = "MTP Scan Day" ;
		SDAY_MTP:actual_range = 20.f, 20.f ;
		SDAY_MTP:Category = "MTP" ;
	float SHOUR_MTP(MTPTime) ;
		SHOUR_MTP:_FillValue = -32767.f ;
		SHOUR_MTP:units = "count" ;
		SHOUR_MTP:long_name = "MTP Scan Hour" ;
		SHOUR_MTP:actual_range = 8.f, 14.f ;
		SHOUR_MTP:Category = "MTP" ;
	float SMIN_MTP(MTPTime) ;
		SMIN_MTP:_FillValue = -32767.f ;
		SMIN_MTP:units = "count" ;
		SMIN_MTP:long_name = "MTP Scan Minute" ;
		SMIN_MTP:actual_range = 0.f, 59.f ;
		SMIN_MTP:Category = "MTP" ;
	float SMONTH_MTP(MTPTime) ;
		SMONTH_MTP:_FillValue = -32767.f ;
		SMONTH_MTP:units = "count" ;
		SMONTH_MTP:long_name = "MTP Scan Month" ;
		SMONTH_MTP:actual_range = 7.f, 7.f ;
		SMONTH_MTP:Category = "MTP" ;
	float SRAT_MTP(MTPTime) ;
		SRAT_MTP:_FillValue = -32767.f ;
		SRAT_MTP:units = "deg_K" ;
		SRAT_MTP:long_name = "MTP Scan RMS Ambient Air Temp" ;
		SRAT_MTP:actual_range = 0.f, 2.01f ;
		SRAT_MTP:Category = "MTP" ;
	float SRLAT_MTP(MTPTime) ;
		SRLAT_MTP:_FillValue = -32767.f ;
		SRLAT_MTP:units = "degree_N" ;
		SRLAT_MTP:long_name = "MTP Scan RMS Latitude" ;
		SRLAT_MTP:actual_range = 0.f, 0.034f ;
		SRLAT_MTP:Category = "MTP" ;
	float SRLON_MTP(MTPTime) ;
		SRLON_MTP:_FillValue = -32767.f ;
		SRLON_MTP:units = "degree_E" ;
		SRLON_MTP:long_name = "MTP Scan RMS Longitude" ;
		SRLON_MTP:actual_range = 0.f, 0.131f ;
		SRLON_MTP:Category = "MTP" ;
	float SRPALT_MTP(MTPTime) ;
		SRPALT_MTP:_FillValue = -32767.f ;
		SRPALT_MTP:units = "km" ;
		SRPALT_MTP:long_name = "MTP Scan RMS Pressure Altitude" ;
		SRPALT_MTP:actual_range = 0.f, 0.08f ;
		SRPALT_MTP:Category = "MTP" ;
	float SRPITCH_MTP(MTPTime) ;
		SRPITCH_MTP:_FillValue = -32767.f ;
		SRPITCH_MTP:units = "degree" ;
		SRPITCH_MTP:long_name = "MTP Scan RMS Pitch" ;
		SRPITCH_MTP:actual_range = 0.01f, 3.08f ;
		SRPITCH_MTP:Category = "MTP" ;
	float SRROLL_MTP(MTPTime) ;
		SRROLL_MTP:_FillValue = -32767.f ;
		SRROLL_MTP:units = "degree" ;
		SRROLL_MTP:long_name = "MTP Scan RMS Roll" ;
		SRROLL_MTP:actual_range = 0.03f, 13.19f ;
		SRROLL_MTP:Category = "MTP" ;
	float SSEC_MTP(MTPTime) ;
		SSEC_MTP:_FillValue = -32767.f ;
		SSEC_MTP:units = "count" ;
		SSEC_MTP:long_name = "MTP Scan Second" ;
		SSEC_MTP:actual_range = 0.f, 59.f ;
		SSEC_MTP:Category = "MTP" ;
	float SYEAR_MTP(MTPTime) ;
		SYEAR_MTP:_FillValue = -32767.f ;
		SYEAR_MTP:units = "count" ;
		SYEAR_MTP:actual_range = 2014.f, 2014.f ;
		SYEAR_MTP:Category = "MTP" ;
///
data:

        CNTSCANANGLE_MTP = 80.f,55.f,42.f,25.f,12.f,0.f,-12.f,-25.f,-42.f,-80.f,-180.f,-180.f ;
	BTSCANANGLE_MTP = 80.f, 55.f,42.f,25.f,12.f,0.f,-12.f,-25.f,-42.f,-80.f ;
        MTPFREQ = 56.363f, 57.612f, 58.363f ;
}
